library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library surf;
use surf.StdRtlPkg.all;

package AesGf2Pkg is

   -- Main operation functionns
   function addRoundKey (state : slv (127 downto 0); key : slv (127 downto 0)) return slv (127 downto 0);
   function subBytes    (state : slv (127 downto 0)) return slv (127 downto 0);
   function shiftRows   (state : slv (127 downto 0)) return slv (127 downto 0);
   function mixColumns  (state : slv (127 downto 0)) return slv (127 downto 0);

   -- Auxialiary functions
   function columnCalculator (column : slv (31 downto 0)) return slv (31 downto 0);
   function subBox           (byte   : slv (7  downto 0)) return slv (7  downto 0);
   function invSubBox        (byte   : slv (7  downto 0)) return slv (7  downto 0);

end AesGf2Pkg;

package body AesGf2Pkg is


   function mixColumns (
      state : slv (127 downto 0)) return slv (127 downto 0) is
      variable output_data : slv (127 downto 0);
   begin
      output_data (31  downto  0) := columnCalculator (state (31  downto  0));
      output_data (63  downto 32) := columnCalculator (state (63  downto 32));
      output_data (95  downto 64) := columnCalculator (state (95  downto 64));
      output_data (127 downto 96) := columnCalculator (state (127 downto 96));
      return output_data;
   end function mixColumns;

   function subBytes (
      state : slv (127 downto 0)) return slv (127 downto 0) is
      variable output_data : slv (127 downto 0);
   begin
      for i 0 to 15 loop
         output_data ((i + 1)*8 - 1 downto i*8) := 
            sBox (state((i + 1)*8 - 1 downto i*8));
      end loop;
      return output_data;
   end function subBytes;

   function shiftRows (
      state : slv (127 downto 0)) return slv (127 downto 0) is
      variable output_data : slv (127 downto 0); 
   begin
      output_data (8*16 - 1 downto 8*15) := state (8*12 - 1 downto 8*11);
      output_data (8*15 - 1 downto 8*14) := state (8*7  - 1 downto  8*6);
      output_data (8*14 - 1 downto 8*13) := state (8*2  - 1 downto  8*1); 
      output_data (8*13 - 1 downto 8*12) := state (8*13 - 1 downto 8*12);
      output_data (8*12 - 1 downto 8*11) := state (8*8  - 1 downto  8*7);
      output_data (8*11 - 1 downto 8*10) := state (8*3  - 1 downto  8*2); 
      output_data (8*10 - 1 downto  8*9) := state (8*14 - 1 downto 8*13);
      output_data (8*9 - 1  downto  8*8) := state (8*9  - 1 downto  8*8);
      output_data (8*8 - 1  downto  8*7) := state (8*4  - 1 downto  8*3);
      output_data (8*7 - 1  downto  8*6) := state (8*15 - 1 downto 8*14);
      output_data (8*6 - 1  downto  8*5) := state (8*10 - 1 downto  8*9);
      output_data (8*5 - 1  downto  8*4) := state (8*5  - 1 downto  8*4);
      output_data (8*4 - 1  downto  8*3) := state (8*16 - 1 downto 8*15);
      output_data (8*3 - 1  downto  8*2) := state (8*11 - 1 downto 8*10);
      output_data (8*2 - 1  downto  8*1) := state (8*6  - 1 downto  8*5);
      output_data (8*1 - 1  downto  8*0) := state (8*1  - 1 downto  8*0); 
      return output_data;
   end function shiftRows;

   function addRoundKey (
      state : slv (127 downto 0);
      key   : slv (127 downto 0)) return slv (127 downto 0) is
   begin
      return state xor key;
   end function addRoundKey;

   function subBox (
      byte : slv (7 downto 0)) return slv (7 downto 0);
   begin
      case byte is
         when x"00" => return x"63";
         when x"01" => return x"7c";
         when x"02" => return x"77";
         when x"03" => return x"7b";
         when x"04" => return x"f2";
         when x"05" => return x"6b";
         when x"06" => return x"6f";
         when x"07" => return x"c5";
         when x"08" => return x"30";
         when x"09" => return x"01";
         when x"0a" => return x"67";
         when x"0b" => return x"2b";
         when x"0c" => return x"fe";
         when x"0d" => return x"d7";
         when x"0e" => return x"ab";
         when x"0f" => return x"76";
         when x"10" => return x"ca";
         when x"11" => return x"82";
         when x"12" => return x"c9";
         when x"13" => return x"7d";
         when x"14" => return x"fa";
         when x"15" => return x"59";
         when x"16" => return x"47";
         when x"17" => return x"f0";
         when x"18" => return x"ad";
         when x"19" => return x"d4";
         when x"1a" => return x"a2";
         when x"1b" => return x"af";
         when x"1c" => return x"9c";
         when x"1d" => return x"a4";
         when x"1e" => return x"72";
         when x"1f" => return x"c0";
         when x"20" => return x"b7";
         when x"21" => return x"fd";
         when x"22" => return x"93";
         when x"23" => return x"26";
         when x"24" => return x"36";
         when x"25" => return x"3f";
         when x"26" => return x"f7";
         when x"27" => return x"cc";
         when x"28" => return x"34";
         when x"29" => return x"a5";
         when x"2a" => return x"e5";
         when x"2b" => return x"f1";
         when x"2c" => return x"71";
         when x"2d" => return x"d8";
         when x"2e" => return x"31";
         when x"2f" => return x"15";
         when x"30" => return x"04";
         when x"31" => return x"c7";
         when x"32" => return x"23";
         when x"33" => return x"c3";
         when x"34" => return x"18";
         when x"35" => return x"96";
         when x"36" => return x"05";
         when x"37" => return x"9a";
         when x"38" => return x"07";
         when x"39" => return x"12";
         when x"3a" => return x"80";
         when x"3b" => return x"e2";
         when x"3c" => return x"eb";
         when x"3d" => return x"27";
         when x"3e" => return x"b2";
         when x"3f" => return x"75";
         when x"40" => return x"09";
         when x"41" => return x"83";
         when x"42" => return x"2c";
         when x"43" => return x"1a";
         when x"44" => return x"1b";
         when x"45" => return x"6e";
         when x"46" => return x"5a";
         when x"47" => return x"a0";
         when x"48" => return x"52";
         when x"49" => return x"3b";
         when x"4a" => return x"d6";
         when x"4b" => return x"b3";
         when x"4c" => return x"29";
         when x"4d" => return x"e3";
         when x"4e" => return x"2f";
         when x"4f" => return x"84";
         when x"50" => return x"53";
         when x"51" => return x"d1";
         when x"52" => return x"00";
         when x"53" => return x"ed";
         when x"54" => return x"20";
         when x"55" => return x"fc";
         when x"56" => return x"b1";
         when x"57" => return x"5b";
         when x"58" => return x"6a";
         when x"59" => return x"cb";
         when x"5a" => return x"be";
         when x"5b" => return x"39";
         when x"5c" => return x"4a";
         when x"5d" => return x"4c";
         when x"5e" => return x"58";
         when x"5f" => return x"cf";
         when x"60" => return x"d0";
         when x"61" => return x"ef";
         when x"62" => return x"aa";
         when x"63" => return x"fb";
         when x"64" => return x"43";
         when x"65" => return x"4d";
         when x"66" => return x"33";
         when x"67" => return x"85";
         when x"68" => return x"45";
         when x"69" => return x"f9";
         when x"6a" => return x"02";
         when x"6b" => return x"7f";
         when x"6c" => return x"50";
         when x"6d" => return x"3c";
         when x"6e" => return x"9f";
         when x"6f" => return x"a8";
         when x"70" => return x"51";
         when x"71" => return x"a3";
         when x"72" => return x"40";
         when x"73" => return x"8f";
         when x"74" => return x"92";
         when x"75" => return x"9d";
         when x"76" => return x"38";
         when x"77" => return x"f5";
         when x"78" => return x"bc";
         when x"79" => return x"b6";
         when x"7a" => return x"da";
         when x"7b" => return x"21";
         when x"7c" => return x"10";
         when x"7d" => return x"ff";
         when x"7e" => return x"f3";
         when x"7f" => return x"d2";
         when x"80" => return x"cd";
         when x"81" => return x"0c";
         when x"82" => return x"13";
         when x"83" => return x"ec";
         when x"84" => return x"5f";
         when x"85" => return x"97";
         when x"86" => return x"44";
         when x"87" => return x"17";
         when x"88" => return x"c4";
         when x"89" => return x"a7";
         when x"8a" => return x"7e";
         when x"8b" => return x"3d";
         when x"8c" => return x"64";
         when x"8d" => return x"5d";
         when x"8e" => return x"19";
         when x"8f" => return x"73";
         when x"90" => return x"60";
         when x"91" => return x"81";
         when x"92" => return x"4f";
         when x"93" => return x"dc";
         when x"94" => return x"22";
         when x"95" => return x"2a";
         when x"96" => return x"90";
         when x"97" => return x"88";
         when x"98" => return x"46";
         when x"99" => return x"ee";
         when x"9a" => return x"b8";
         when x"9b" => return x"14";
         when x"9c" => return x"de";
         when x"9d" => return x"5e";
         when x"9e" => return x"0b";
         when x"9f" => return x"db";
         when x"a0" => return x"e0";
         when x"a1" => return x"32";
         when x"a2" => return x"3a";
         when x"a3" => return x"0a";
         when x"a4" => return x"49";
         when x"a5" => return x"06";
         when x"a6" => return x"24";
         when x"a7" => return x"5c";
         when x"a8" => return x"c2";
         when x"a9" => return x"d3";
         when x"aa" => return x"ac";
         when x"ab" => return x"62";
         when x"ac" => return x"91";
         when x"ad" => return x"95";
         when x"ae" => return x"e4";
         when x"af" => return x"79";
         when x"b0" => return x"e7";
         when x"b1" => return x"c8";
         when x"b2" => return x"37";
         when x"b3" => return x"6d";
         when x"b4" => return x"8d";
         when x"b5" => return x"d5";
         when x"b6" => return x"4e";
         when x"b7" => return x"a9";
         when x"b8" => return x"6c";
         when x"b9" => return x"56";
         when x"ba" => return x"f4";
         when x"bb" => return x"ea";
         when x"bc" => return x"65";
         when x"bd" => return x"7a";
         when x"be" => return x"ae";
         when x"bf" => return x"08";
         when x"c0" => return x"ba";
         when x"c1" => return x"78";
         when x"c2" => return x"25";
         when x"c3" => return x"2e";
         when x"c4" => return x"1c";
         when x"c5" => return x"a6";
         when x"c6" => return x"b4";
         when x"c7" => return x"c6";
         when x"c8" => return x"e8";
         when x"c9" => return x"dd";
         when x"ca" => return x"74";
         when x"cb" => return x"1f";
         when x"cc" => return x"4b";
         when x"cd" => return x"bd";
         when x"ce" => return x"8b";
         when x"cf" => return x"8a";
         when x"d0" => return x"70";
         when x"d1" => return x"3e";
         when x"d2" => return x"b5";
         when x"d3" => return x"66";
         when x"d4" => return x"48";
         when x"d5" => return x"03";
         when x"d6" => return x"f6";
         when x"d7" => return x"0e";
         when x"d8" => return x"61";
         when x"d9" => return x"35";
         when x"da" => return x"57";
         when x"db" => return x"b9";
         when x"dc" => return x"86";
         when x"dd" => return x"c1";
         when x"de" => return x"1d";
         when x"df" => return x"9e";
         when x"e0" => return x"e1";
         when x"e1" => return x"f8";
         when x"e2" => return x"98";
         when x"e3" => return x"11";
         when x"e4" => return x"69";
         when x"e5" => return x"d9";
         when x"e6" => return x"8e";
         when x"e7" => return x"94";
         when x"e8" => return x"9b";
         when x"e9" => return x"1e";
         when x"ea" => return x"87";
         when x"eb" => return x"e9";
         when x"ec" => return x"ce";
         when x"ed" => return x"55";
         when x"ee" => return x"28";
         when x"ef" => return x"df";
         when x"f0" => return x"8c";
         when x"f1" => return x"a1";
         when x"f2" => return x"89";
         when x"f3" => return x"0d";
         when x"f4" => return x"bf";
         when x"f5" => return x"e6";
         when x"f6" => return x"42";
         when x"f7" => return x"68";
         when x"f8" => return x"41";
         when x"f9" => return x"99";
         when x"fa" => return x"2d";
         when x"fb" => return x"0f";
         when x"fc" => return x"b0";
         when x"fd" => return x"54";
         when x"fe" => return x"bb";
         when x"ff" => return x"16";
         when others => return (others => '0');
      end case;
   end function subBox;

   function invSubBox(
      byte : slv(7 downto 0)) return slv is
   begin
      case byte is
         when x"00" => return x"52";
         when x"01" => return x"09";
         when x"02" => return x"6A";
         when x"03" => return x"D5";
         when x"04" => return x"30";
         when x"05" => return x"36";
         when x"06" => return x"A5";
         when x"07" => return x"38";
         when x"08" => return x"BF";
         when x"09" => return x"40";
         when x"0A" => return x"A3";
         when x"0B" => return x"9E";
         when x"0C" => return x"81";
         when x"0D" => return x"F3";
         when x"0E" => return x"D7";
         when x"0F" => return x"FB";
         when x"10" => return x"7C";
         when x"11" => return x"E3";
         when x"12" => return x"39";
         when x"13" => return x"82";
         when x"14" => return x"9B";
         when x"15" => return x"2F";
         when x"16" => return x"FF";
         when x"17" => return x"87";
         when x"18" => return x"34";
         when x"19" => return x"8E";
         when x"1A" => return x"43";
         when x"1B" => return x"44";
         when x"1C" => return x"C4";
         when x"1D" => return x"DE";
         when x"1E" => return x"E9";
         when x"1F" => return x"CB";
         when x"20" => return x"54";
         when x"21" => return x"7B";
         when x"22" => return x"94";
         when x"23" => return x"32";
         when x"24" => return x"A6";
         when x"25" => return x"C2";
         when x"26" => return x"23";
         when x"27" => return x"3D";
         when x"28" => return x"EE";
         when x"29" => return x"4C";
         when x"2A" => return x"95";
         when x"2B" => return x"0B";
         when x"2C" => return x"42";
         when x"2D" => return x"FA";
         when x"2E" => return x"C3";
         when x"2F" => return x"4E";
         when x"30" => return x"08";
         when x"31" => return x"2E";
         when x"32" => return x"A1";
         when x"33" => return x"66";
         when x"34" => return x"28";
         when x"35" => return x"D9";
         when x"36" => return x"24";
         when x"37" => return x"B2";
         when x"38" => return x"76";
         when x"39" => return x"5B";
         when x"3A" => return x"A2";
         when x"3B" => return x"49";
         when x"3C" => return x"6D";
         when x"3D" => return x"8B";
         when x"3E" => return x"D1";
         when x"3F" => return x"25";
         when x"40" => return x"72";
         when x"41" => return x"F8";
         when x"42" => return x"F6";
         when x"43" => return x"64";
         when x"44" => return x"86";
         when x"45" => return x"68";
         when x"46" => return x"98";
         when x"47" => return x"16";
         when x"48" => return x"D4";
         when x"49" => return x"A4";
         when x"4A" => return x"5C";
         when x"4B" => return x"CC";
         when x"4C" => return x"5D";
         when x"4D" => return x"65";
         when x"4E" => return x"B6";
         when x"4F" => return x"92";
         when x"50" => return x"6C";
         when x"51" => return x"70";
         when x"52" => return x"48";
         when x"53" => return x"50";
         when x"54" => return x"FD";
         when x"55" => return x"ED";
         when x"56" => return x"B9";
         when x"57" => return x"DA";
         when x"58" => return x"5E";
         when x"59" => return x"15";
         when x"5A" => return x"46";
         when x"5B" => return x"57";
         when x"5C" => return x"A7";
         when x"5D" => return x"8D";
         when x"5E" => return x"9D";
         when x"5F" => return x"84";
         when x"60" => return x"90";
         when x"61" => return x"D8";
         when x"62" => return x"AB";
         when x"63" => return x"00";
         when x"64" => return x"8C";
         when x"65" => return x"BC";
         when x"66" => return x"D3";
         when x"67" => return x"0A";
         when x"68" => return x"F7";
         when x"69" => return x"E4";
         when x"6A" => return x"58";
         when x"6B" => return x"05";
         when x"6C" => return x"B8";
         when x"6D" => return x"B3";
         when x"6E" => return x"45";
         when x"6F" => return x"06";
         when x"70" => return x"D0";
         when x"71" => return x"2C";
         when x"72" => return x"1E";
         when x"73" => return x"8F";
         when x"74" => return x"CA";
         when x"75" => return x"3F";
         when x"76" => return x"0F";
         when x"77" => return x"02";
         when x"78" => return x"C1";
         when x"79" => return x"AF";
         when x"7A" => return x"BD";
         when x"7B" => return x"03";
         when x"7C" => return x"01";
         when x"7D" => return x"13";
         when x"7E" => return x"8A";
         when x"7F" => return x"6B";
         when x"80" => return x"3A";
         when x"81" => return x"91";
         when x"82" => return x"11";
         when x"83" => return x"41";
         when x"84" => return x"4F";
         when x"85" => return x"67";
         when x"86" => return x"DC";
         when x"87" => return x"EA";
         when x"88" => return x"97";
         when x"89" => return x"F2";
         when x"8A" => return x"CF";
         when x"8B" => return x"CE";
         when x"8C" => return x"F0";
         when x"8D" => return x"B4";
         when x"8E" => return x"E6";
         when x"8F" => return x"73";
         when x"90" => return x"96";
         when x"91" => return x"AC";
         when x"92" => return x"74";
         when x"93" => return x"22";
         when x"94" => return x"E7";
         when x"95" => return x"AD";
         when x"96" => return x"35";
         when x"97" => return x"85";
         when x"98" => return x"E2";
         when x"99" => return x"F9";
         when x"9A" => return x"37";
         when x"9B" => return x"E8";
         when x"9C" => return x"1C";
         when x"9D" => return x"75";
         when x"9E" => return x"DF";
         when x"9F" => return x"6E";
         when x"A0" => return x"47";
         when x"A1" => return x"F1";
         when x"A2" => return x"1A";
         when x"A3" => return x"71";
         when x"A4" => return x"1D";
         when x"A5" => return x"29";
         when x"A6" => return x"C5";
         when x"A7" => return x"89";
         when x"A8" => return x"6F";
         when x"A9" => return x"B7";
         when x"AA" => return x"62";
         when x"AB" => return x"0E";
         when x"AC" => return x"AA";
         when x"AD" => return x"18";
         when x"AE" => return x"BE";
         when x"AF" => return x"1B";
         when x"B0" => return x"FC";
         when x"B1" => return x"56";
         when x"B2" => return x"3E";
         when x"B3" => return x"4B";
         when x"B4" => return x"C6";
         when x"B5" => return x"D2";
         when x"B6" => return x"79";
         when x"B7" => return x"20";
         when x"B8" => return x"9A";
         when x"B9" => return x"DB";
         when x"BA" => return x"C0";
         when x"BB" => return x"FE";
         when x"BC" => return x"78";
         when x"BD" => return x"CD";
         when x"BE" => return x"5A";
         when x"BF" => return x"F4";
         when x"C0" => return x"1F";
         when x"C1" => return x"DD";
         when x"C2" => return x"A8";
         when x"C3" => return x"33";
         when x"C4" => return x"88";
         when x"C5" => return x"07";
         when x"C6" => return x"C7";
         when x"C7" => return x"31";
         when x"C8" => return x"B1";
         when x"C9" => return x"12";
         when x"CA" => return x"10";
         when x"CB" => return x"59";
         when x"CC" => return x"27";
         when x"CD" => return x"80";
         when x"CE" => return x"EC";
         when x"CF" => return x"5F";
         when x"D0" => return x"60";
         when x"D1" => return x"51";
         when x"D2" => return x"7F";
         when x"D3" => return x"A9";
         when x"D4" => return x"19";
         when x"D5" => return x"B5";
         when x"D6" => return x"4A";
         when x"D7" => return x"0D";
         when x"D8" => return x"2D";
         when x"D9" => return x"E5";
         when x"DA" => return x"7A";
         when x"DB" => return x"9F";
         when x"DC" => return x"93";
         when x"DD" => return x"C9";
         when x"DE" => return x"9C";
         when x"DF" => return x"EF";
         when x"E0" => return x"A0";
         when x"E1" => return x"E0";
         when x"E2" => return x"3B";
         when x"E3" => return x"4D";
         when x"E4" => return x"AE";
         when x"E5" => return x"2A";
         when x"E6" => return x"F5";
         when x"E7" => return x"B0";
         when x"E8" => return x"C8";
         when x"E9" => return x"EB";
         when x"EA" => return x"BB";
         when x"EB" => return x"3C";
         when x"EC" => return x"83";
         when x"ED" => return x"53";
         when x"EE" => return x"99";
         when x"EF" => return x"61";
         when x"F0" => return x"17";
         when x"F1" => return x"2B";
         when x"F2" => return x"04";
         when x"F3" => return x"7E";
         when x"F4" => return x"BA";
         when x"F5" => return x"77";
         when x"F6" => return x"D6";
         when x"F7" => return x"26";
         when x"F8" => return x"E1";
         when x"F9" => return x"69";
         when x"FA" => return x"14";
         when x"FB" => return x"63";
         when x"FC" => return x"55";
         when x"FD" => return x"21";
         when x"FE" => return x"0C";
         when x"FF" => return x"7D";
         when others => return (others => '0');
      end case;
   end function invSubBox;

end package body AesGf2Pkg;
